`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06.05.2022 07:46:06
// Design Name: 
// Module Name: Display7
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Display7(
    input CLK,
    input [3:0] ADC,
    output reg [13:0] D7);
    
    always @(*)
        case(ADC)
            4'b0000: D7=14'b00000010000001;//0
            4'b0001: D7=14'b00000011001111;//1
            4'b0010: D7=14'b00000010010010;//2
            4'b0011: D7=14'b00000010000110;//3
            4'b0100: D7=14'b00000011001100;//4
            4'b0101: D7=14'b00000010100100;//5
            4'b0110: D7=14'b00000010100000;//6
            4'b0111: D7=14'b00000010001111;//7
            4'b1000: D7=14'b00000010000000;//8
            4'b1001: D7=14'b00000010000100;//9
            4'b1010: D7=14'b10011110000001;//10
            4'b1011: D7=14'b10011111001111;//11
            4'b1100: D7=14'b10011110010010;//12
            4'b1101: D7=14'b10011110000110;//13
            4'b1110: D7=14'b10011111001100;//14
            4'b1111: D7=14'b10011110100100;//15
        endcase
endmodule
